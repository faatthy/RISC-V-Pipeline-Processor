module ADDER(
    input [31:0]A,B,
    output  [31:0]y
);
assign y=A+B;
endmodule
